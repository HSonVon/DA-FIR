module top_SDA (
    input CLOCK_50,
    input [0:0] KEY,
    output signed [15:0] Yn
);
    reg signed [7:0] X;    
    reg [7:0] addr;
    reg [3:0] delay_counter;
    reg delayed_output;

    SDA8FIR sdafir (
        .clk(CLOCK_50),
        .RstN(KEY[0:0]),
        .X(X),
        .Yn(Yn)
    );

    always @(posedge CLOCK_50 or negedge KEY[0:0]) begin
        if (!KEY[0:0]) begin
            addr = 8'd0;
            delay_counter = 4'd0;
            delayed_output = 1'b0;
        end else begin
            if (delay_counter < 4'd8) begin
                delay_counter = delay_counter + 4'd1;
            end else begin
                delay_counter = 4'd0;
                delayed_output = 1'b1;
                addr = (addr == 8'd176) ? 8'd0 : addr + 8'd1;
            end
        end
    end

    always @(*) begin
        if (!KEY[0:0]) begin
            X = 8'd0;
        end else if (delayed_output) begin
            case (addr)
                8'd0: X = 8'd0;
                8'd1: X = 8'd127;
                8'd2: X = 8'd107;
                8'd3: X = -8'd28;
                8'd4: X = -8'd60;
                8'd5: X = 8'd75;
                8'd6: X = 8'd127;
                8'd7: X = 8'd127;
                8'd8: X = 8'd33;
                8'd9: X = -8'd6;
                8'd10: X = 8'd122;
                8'd11: X = 8'd127;
                8'd12: X = 8'd127;
                8'd13: X = 8'd53;
                8'd14: X = 8'd4;
                8'd15: X = 8'd122;
                8'd16: X = 8'd127;
                8'd17: X = 8'd127;
                8'd18: X = 8'd23;
                8'd19: X = -8'd34;
                8'd20: X = 8'd75;
                8'd21: X = 8'd127;
                8'd22: X = 8'd122;
                8'd23: X = -8'd43;
                8'd24: X = -8'd106;
                8'd25: X = 8'd0;
                8'd26: X = 8'd106;
                8'd27: X = 8'd43;
                8'd28: X = -8'd122;
                8'd29: X = -8'd128;
                8'd30: X = -8'd75;
                8'd31: X = 8'd34;
                8'd32: X = -8'd23;
                8'd33: X = -8'd128;
                8'd34: X = -8'd128;
                8'd35: X = -8'd122;
                8'd36: X = -8'd4;
                8'd37: X = -8'd53;
                8'd38: X = -8'd128;
                8'd39: X = -8'd128;
                8'd40: X = -8'd122;
                8'd41: X = 8'd6;
                8'd42: X = -8'd33;
                8'd43: X = -8'd128;
                8'd44: X = -8'd128;
                8'd45: X = -8'd75;
                8'd46: X = 8'd60;
                8'd47: X = 8'd28;
                8'd48: X = -8'd107;
                8'd49: X = -8'd128;
                8'd50: X = 8'd0;
                8'd51: X = 8'd127;
                8'd52: X = 8'd107;
                8'd53: X = -8'd28;
                8'd54: X = -8'd60;
                8'd55: X = 8'd75;
                8'd56: X = 8'd127;
                8'd57: X = 8'd127;
                8'd58: X = 8'd33;
                8'd59: X = -8'd6;
                8'd60: X = 8'd122;
                8'd61: X = 8'd127;
                8'd62: X = 8'd127;
                8'd63: X = 8'd53;
                8'd64: X = 8'd4;
                8'd65: X = 8'd122;
                8'd66: X = 8'd127;
                8'd67: X = 8'd127;
                8'd68: X = 8'd23;
                8'd69: X = -8'd34;
                8'd70: X = 8'd75;
                8'd71: X = 8'd127;
                8'd72: X = 8'd122;
                8'd73: X = -8'd43;
                8'd74: X = -8'd106;
                8'd75: X = 8'd0;
                8'd76: X = 8'd106;
                8'd77: X = 8'd43;
                8'd78: X = -8'd122;
                8'd79: X = -8'd128;
                8'd80: X = -8'd75;
                8'd81: X = 8'd34;
                8'd82: X = -8'd23;
                8'd83: X = -8'd128;
                8'd84: X = -8'd128;
                8'd85: X = -8'd122;
                8'd86: X = -8'd4;
                8'd87: X = -8'd53;
                8'd88: X = -8'd128;
                8'd89: X = -8'd128;
                8'd90: X = -8'd122;
                8'd91: X = 8'd6;
                8'd92: X = -8'd33;
                8'd93: X = -8'd128;
                8'd94: X = -8'd128;
                8'd95: X = -8'd75;
                8'd96: X = 8'd60;
                8'd97: X = 8'd28;
                8'd98: X = -8'd107;
                8'd99: X = -8'd128;
                8'd100: X = 8'd0;
                8'd101: X = 8'd127;
                8'd102: X = 8'd107;
                8'd103: X = -8'd28;
                8'd104: X = -8'd60;
                8'd105: X = 8'd75;
                8'd106: X = 8'd127;
                8'd107: X = 8'd127;
                8'd108: X = 8'd33;
                8'd109: X = -8'd6;
                8'd110: X = 8'd122;
                8'd111: X = 8'd127;
                8'd112: X = 8'd127;
                8'd113: X = 8'd53;
                8'd114: X = 8'd4;
                8'd115: X = 8'd122;
                8'd116: X = 8'd127;
                8'd117: X = 8'd127;
                8'd118: X = 8'd23;
                8'd119: X = -8'd34;
                8'd120: X = 8'd75;
                8'd121: X = 8'd127;
                8'd122: X = 8'd122;
                8'd123: X = -8'd43;
                8'd124: X = -8'd106;
                8'd125: X = 8'd0;
                8'd126: X = 8'd106;
                8'd127: X = 8'd43;
                8'd128: X = -8'd122;
                8'd129: X = -8'd128;
                8'd130: X = -8'd75;
                8'd131: X = 8'd34;
                8'd132: X = -8'd23;
                8'd133: X = -8'd128;
                8'd134: X = -8'd128;
                8'd135: X = -8'd122;
                8'd136: X = -8'd4;
                8'd137: X = -8'd53;
                8'd138: X = -8'd128;
                8'd139: X = -8'd128;
                8'd140: X = -8'd122;
                8'd141: X = 8'd6;
                8'd142: X = -8'd33;
                8'd143: X = -8'd128;
                8'd144: X = -8'd128;
                8'd145: X = -8'd75;
                8'd146: X = 8'd60;
                8'd147: X = 8'd28;
                8'd148: X = -8'd107;
                8'd149: X = -8'd128;
                8'd150: X = 8'd0;
                8'd151: X = 8'd127;
                8'd152: X = 8'd107;
                8'd153: X = -8'd28;
                8'd154: X = -8'd60;
                8'd155: X = 8'd75;
                8'd156: X = 8'd127;
                8'd157: X = 8'd127;
                8'd158: X = 8'd33;
                8'd159: X = -8'd6;
                8'd160: X = 8'd122;
                8'd161: X = 8'd127;
                8'd162: X = 8'd127;
                8'd163: X = 8'd53;
                8'd164: X = 8'd4;
                8'd165: X = 8'd122;
                8'd166: X = 8'd127;
                8'd167: X = 8'd127;
                8'd168: X = 8'd23;
                8'd169: X = -8'd34;
                8'd170: X = 8'd75;
                8'd171: X = 8'd127;
                8'd172: X = 8'd122;
                8'd173: X = -8'd43;
                8'd174: X = -8'd106;
                8'd175: X = 8'd0;
                8'd176: X = 8'd106;
                default: X = 8'd0;
            endcase
        end
    end
endmodule 